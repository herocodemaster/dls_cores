
/* verilator lint_restore */
/* verilator tracing_on */
/* verilator coverage_on */

