
module dlsc_empty;

endmodule

