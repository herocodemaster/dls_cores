// 
// Copyright (c) 2011, Daniel Strother < http://danstrother.com/ >
// All rights reserved.
// 
// Redistribution and use in source and binary forms, with or without
// modification, are permitted provided that the following conditions are met:
//   - Redistributions of source code must retain the above copyright notice,
//     this list of conditions and the following disclaimer.
//   - Redistributions in binary form must reproduce the above copyright
//     notice, this list of conditions and the following disclaimer in the
//     documentation and/or other materials provided with the distribution.
//   - The name of the author may not be used to endorse or promote products
//     derived from this software without specific prior written permission.
// 
// THIS SOFTWARE IS PROVIDED BY THE AUTHOR "AS IS" AND ANY EXPRESS OR IMPLIED
// WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED WARRANTIES OF
// MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE DISCLAIMED. IN NO
// EVENT SHALL THE AUTHOR BE LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL,
// SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED
// TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES; LOSS OF USE, DATA, OR
// PROFITS; OR BUSINESS INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF
// LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT (INCLUDING
// NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE OF THIS
// SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
//


// some tools support $clog2, but don't support constant functions (Icarus and Covered)
// other tools support constant functions, but don't support $clog2 (XST)
// ..hence the `ifdef
`ifdef USE_CLOG2

    `define dlsc_clog2(x) $clog2(x)

    `define dlsc_clog2_lower(x,lower_bound) (($clog2(x) < (lower_bound)) ? (lower_bound) : $clog2(x))
    `define dlsc_clog2_upper(x,upper_bound) (($clog2(x) > (upper_bound)) ? (upper_bound) : $clog2(x))

`else

    `define dlsc_clog2(x) dlsc_clog2_func(x)
    
    `define dlsc_clog2_lower(x,lower_bound) ((dlsc_clog2_func(x) < (lower_bound)) ? (lower_bound) : dlsc_clog2_func(x))
    `define dlsc_clog2_upper(x,upper_bound) ((dlsc_clog2_func(x) > (upper_bound)) ? (upper_bound) : dlsc_clog2_func(x))

    function integer dlsc_clog2_func;
        input integer val;
        integer i;
    begin
        i = val - 1;
        for(dlsc_clog2_func=0;i>0;dlsc_clog2_func=dlsc_clog2_func+1)
            i = i >> 1;
    end
    endfunction

`endif

