
/* verilator coverage_off */
/* verilator tracing_off */
/* verilator lint_off WIDTH */
`include "dlsc_sim.vh"

