
/* verilator lint_on WIDTH */
/* verilator tracing_on */
/* verilator coverage_on */

