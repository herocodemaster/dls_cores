
/* verilator coverage_off */
/* verilator tracing_off */
/* verilator lint_save */
/* verilator lint_off WIDTH */
/* verilator lint_off BLKSEQ */
/* verilator lint_off UNUSED */
`include "dlsc_sim.vh"

